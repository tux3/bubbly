`default_nettype none

