`include "core/params.svh"

// Location of the boot code in flash (4MiB)
`define FLASH_TEXT_ADDR 'h400000

module top(
    input CLK100MHZ,
    input RSTN,

    // SPI_CLK is on a non-CCIO pin, it can't be routed to a BUFG...
    (* clock_buffer_type = "BUFR" *)
    input SPI_CLK,
    input SPI_MOSI,
    output SPI_MISO,
    input SPI_SS,

    output FLASH_CS,
    output FLASH_CLK,
    inout FLASH_MOSI,
    inout FLASH_MISO,
    inout FLASH_WP,
    inout FLASH_HOLD,
    
    input ETH_COL,
    input ETH_CRS,
    output ETH_REF_CLK,
    output ETH_RSTN,
    input ETH_RX_CLK,
    input ETH_RX_DV,
    input [3:0] ETH_RXD,
    input ETH_RXERR,
    input ETH_TX_CLK,
    output ETH_TX_EN,
    output [3:0] ETH_TXD,

    input [3:0] SWITCH,
    output [9:0] PROBE,
    output PROBE_GND_34,
    output reg [3:0] LED
    );

wire clk, rst;
wire flash_capture_clk;
wire eth_ref_clk;
assign ETH_REF_CLK = eth_ref_clk;
pll pll(
    .CLK100MHZ,
    .RSTN,
    .clk,
    .rst,
    .flash_capture_clk,
    .eth_ref_clk
);

reg [$bits(SWITCH)-1:0] switch_sync1;
reg [$bits(SWITCH)-1:0] switch_reg;
always_ff @(posedge flash_capture_clk) begin
    switch_sync1 <= SWITCH;
    switch_reg <= switch_sync1;
end

spi_soc #(.RESET_PC(`FLASH_TEXT_ADDR)) spi_soc(
    .clk,
    .rst,
    
    .ETH_RX_CLK(ETH_RX_CLK),
    .ETH_RXD(ETH_RXD),
    .ETH_RX_DV(ETH_RX_DV),
    .ETH_RXERR(ETH_RXERR),
    .ETH_TX_CLK(ETH_TX_CLK),
    .ETH_TXD(ETH_TXD),
    .ETH_TX_EN(ETH_TX_EN),
    .ETH_COL(ETH_COL),
    .ETH_CRS(ETH_CRS),
    .ETH_RSTN(ETH_RSTN),

    .FLASH_CAPTURE_CLK(flash_capture_clk),

    .SWITCH(switch_reg[0]),
    .PROBE,
    .LED(LED[3:1]),

    .*
);

assign PROBE_GND_34 = '0;

logic [24:0] counter;
assign LED[0] = counter[$bits(counter)-1];

always_ff @(posedge clk) begin
    if (rst)
        counter <= '0;
    else
        counter <= counter + 1;
end

endmodule
